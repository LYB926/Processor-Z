//存储器文件ram.v
module ram(
input               clock,
input[8:0]          addr,
input               wr,
input[31:0]         wdata,
input               rd,
output reg[31:0]    rdata
);
//TBD

endmodule