//寄存器读写文件 regfile.v
module regfile(
input[3:0]      dstE,
input[31:0]     valE,
input[3:0]      dstM,
input[31:0]     valM,
input           reset,
input           clock,
output[31:0]    r0,
output[31:0]    r1,
output[31:0]    r2,
output[31:0]    r3,
output[31:0]    r4,
output[31:0]    r5,
output[31:0]    r6,
output[31:0]    r7
);
//TBD

endmodule